///////////////////////////////////////////////
//Company: ITESO
//Engineer: Antonio Rangel Avila  
//Module Description: Data path, RISC-V 32bits multi-cycle,parameterized;
//Date: March 4th 2023
///////////////////////////////////////////////
module Data_Path #(parameter DATA_WIDTH = 32)(
//INPUTS
input clk, reset,

//CONTROL SIGNALS
input IRWrite, 			//The instruction code is stored here
input [3:0] ALUControl, //Add base address to offset
input IorD,					//Load data from memory
input RegWrite,         //Write Data to register file
input [1:0] ALUSrcA,    //Increment PC by 4 or 1 
input [1:0] ALUSrcB,    //Increment PC by 4 or 1
input MemWrite,         //Enhanced datapath for sw instruction
//input [1:0]RegDst,    //Enhanced datapath for R-type instruction
input [1:0] MemtoReg,   //Enhanced datapath for R-type instruction
input PCEn,					//enhanced for beq instruction
input [1:0] PCSrc,   	//enhanced for beq instruction

output Zero,
output [6:0] Op,
output [2:0] Funct3,
output [6:0] Funct7,

input [7:0] gpio_port_in,   //GPIO Ports
output [7:0] gpio_port_out, //GPIO Ports

input uart_rx, 				//UART Ports
output uart_tx 				//UART Ports

);

wire [DATA_WIDTH-1:0] pc, pc_next;
wire [DATA_WIDTH-1:0] ALUOut;
wire [DATA_WIDTH-1:0] Adr;
wire [DATA_WIDTH-1:0] Read_Data;

wire [DATA_WIDTH-1:0] Instr;

//-----New wires added for risc-v-32I implementation
wire [6:0] op_d, op_q;
wire [2:0] funct3_d, funct3_q;
wire [6:0] funct7_d, funct7_q;
wire [4:0] rs1_d, rs1_q;
wire [4:0] rs2_d, rs2_q;
wire [4:0] rd_d, rd_q;
wire [11:0] imm_d, imm_q;
//-----could be no used:
/*wire [3:0] shamt;
wire [6:0] csr;
wire branch;
wire jal;
wire jalr;
wire load;
wire store;
wire alu;
wire [1:0] mem_size;
wire [1:0] mem_signed;*/

 
//--------------------------------------------------
wire [DATA_WIDTH-1:0] Write_Data;
//wire [4:0] Write_Register;
wire [DATA_WIDTH-1:0] Data;
wire [DATA_WIDTH-1:0] rd1, rd2, a, b;
wire [DATA_WIDTH-1:0] SrcA, SrcB;
wire [DATA_WIDTH-1:0] ALUResult;
wire [DATA_WIDTH-1:0] Sign_Imm;
wire [DATA_WIDTH-1:0] Shifted_Imm;
wire [DATA_WIDTH-1:0] OldPC;
//--------------------------------------------------
wire RAMen, GPIOen, UARTen;
wire [DATA_WIDTH-1:0] NADDR, FromMem, GPIOData, ROMDataOut, ram_out, UARTData;
wire [1:0] DataSel;
//--------------------------------------------------
Reg_param  #
					(

								 .reset_value(32'h400000)
					) 
					Pc 
					(
								 .rst(reset), 
								 .clk(clk), 
								 .enable(PCEn), 
								 .D(pc_next), 
								 .Q(pc)
					);
					
Mux2x1 instr_or_data (
								 .Selector(IorD),
								 .I_0(pc),
								 .I_1(ALUOut),
								 .Mux_Out(Adr)
						   );
							
Memory_Controller #
					(
								.DATA_WIDTH(32), .ADDR_WIDTH(32)
					) 
					MemCtrl
					(
								.WrtEn(MemWrite),
								.ADDRIn(Adr),
								.RAM_En(RAMen),
								.GPIO_En(GPIOen),
								.UART_En(UARTen),
								.Sel(DataSel),
								.ADDROut(NADDR)
					);
					
Mux4x1 peripheral_mux ( 
								.Selector(DataSel), 
								.I_0(ram_out), 
								.I_1(UARTData), 
								.I_2(GPIOData), 
								.I_3(ROMDataOut), 
								.Mux_Out(Read_Data)
							);
					
Data_Memory		RAM 	(
								.clk				(clk),
								.Write_Enable	(RAMen),
								.Write_Data		(b),						
								.Address       (NADDR),
								.Read_Data		(ram_out)
							);
UART uart_0
							(
								.clk(clk),
								.rst(reset),
								.wrtEn(UARTen),
								.addr(NADDR[2]),
								.TxData(b),
								.ReadReg(UARTData),
								.SerialOut(uart_tx),
								.SerialIn(uart_rx)
							);
							
GPIO gpio_0				(
								.clk(clk),
								.rst(reset),
								.en(GPIOen),
								.addr(NADDR[2]), 
								.PORT_IN(gpio_port_in),
								.DataToOut(b),
								.PORT_OUT(gpio_port_out),
								.DataFromIn(GPIOData)
							);
							
Program_Memory	ROM	(
									.Address			(NADDR),
									.Instruction	(ROMDataOut)
								);

							
/*Memory_System ROM_RAM (
                         .clk(clk),
								 .Write_Enable_i(MemWrite),
								 .Write_Data_i(b),
								 .Address_i(Adr),
								 .Instruction_o(Read_Data)
                      ); */
							 
Decoder Decoder_rv32I (
								 .instr(Read_Data), //input
								 
								 .opcode(op_d),
								 .funct3(funct3_d),
								 .funct7(funct7_d),
								 .rs1(rs1_d),
								 .rs2(rs2_d),
								 .rd(rd_d),
								 .imm(imm_d)
								 /*.shamt(),
								 .csr(),
								 .branch(),
								 .jal(),
								 .jalr(),
								 .load(),
								 .store(),
								 .alu(),
								 .mem_size(),
								 .mem_signed()*/

                      );
							 

			

Reg_param #(.width(7)) IR_opcode (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite),	
																			.D(op_d),	
																			.Q(op_q)
																	  );
																	  
Reg_param #(.width(5)) IR_rd (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite),	
																			.D(rd_d),	
																			.Q(rd_q)
																	  );
																	  
Reg_param #(.width(5)) IR_rs1 (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite),	
																			.D(rs1_d),	
																			.Q(rs1_q)
																	  );
																	  
Reg_param #(.width(5)) IR_rs2 (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite),	
																			.D(rs2_d),	
																			.Q(rs2_q)
																	  );
																	  
Reg_param #(.width(3)) IR_funct3 (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite),	
																			.D(funct3_d),	
																			.Q(funct3_q)
																	  );
Reg_param #(.width(7)) IR_funct7 (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite),	
																			.D(funct7_d),	
																			.Q(funct7_q)
																	  );
																	  
Reg_param #(.width(12)) IR_imm (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite),	
																			.D(imm_d),	
																			.Q(imm_q)
																	  );
																	  
Reg_param old_PC (
																			.rst(reset), 
																			.clk(clk), 
																			.enable(IRWrite), 
																			.D(pc), 
																			.Q(OldPC)
																	  );
													
																	  
																	  

Reg_param Memory_Data_register (
											.rst(reset), 
											.clk(clk), 
											.enable(1'b1), 
											.D(Read_Data), 
											.Q(Data)
								);
								 
/*Mux4x1  #(.DATA_WIDTH(5)) Rrt_or_Rrd (
													.Selector(RegDst), 
													.I_0(Instr[20:16]), 
													.I_1(Instr[15:11]), 
													.I_2(5'd31), 
													.I_3(5'd0), 
													.Mux_Out(Write_Register)
												 );*/

Mux4x1 Write_data_mux ( 
													.Selector(MemtoReg), 
													.I_0(ALUOut), 
													.I_1(Data), 
													.I_2(32'b0), 
													.I_3(32'b0), 
													.Mux_Out(Write_Data)
						    );
							 
rv32i_imm_gen imm_gen  (
												  .opcode(op_q),
												  .funct3(funct3_q),
												  .rs1(rs1_q),
												  .rs2(rs2_q),
												  .rd(rd_q),
												  .funct7(funct7_q),
												  .imm_in(imm_q),
												  .imm(Sign_Imm)
												);
								
							
Reg_File Reg_file (
													.A1(rs1_q),  
													.A2(rs2_q), 
													.A3(rd_q),
												   .rst(reset), .clk(clk), 
											   	.WE3(RegWrite), .WD3(Write_Data),
													.RD1(rd1), .RD2(rd2)
                  );
						
Reg_param A_Register (
													.rst(reset), 
													.clk(clk), 
													.enable(1'b1), 
													.D(rd1), 
													.Q(a)
							);
							
Reg_param B_Register (
													.rst(reset), 
													.clk(clk), 
													.enable(1'b1), 
													.D(rd2), 
													.Q(b)
							);
							
/*Sign_Extend	Sign_Ext	(
									.Imm				(Instr[15:0]),
									.Sign_Ext_Imm	(Sign_Imm)
							);
	
Shift_Left_2 Branch_Shift	(
											.Ext_Imm			(Sign_Imm),
											.Shifted_Imm	(Shifted_Imm)
									);*/
							
/*Mux2x1 mux_a_input   (
								 .Selector(ALUSrcA),
								 .I_0(pc),
								 .I_1(a),
								 .Mux_Out(SrcA)
						   ); */
							
Mux4x1 mux_a_input    ( 
													.Selector(ALUSrcA), 
													.I_0(pc), 
													.I_1(a), 
													.I_2(OldPC), 
													.I_3(32'h0), 
													.Mux_Out(SrcA)
						    );							
							
Mux4x1 mux_b_input    ( 
													.Selector(ALUSrcB), 
													.I_0(b), 
													.I_1(4), 
													.I_2(Sign_Imm), 
													.I_3(0), 
													.Mux_Out(SrcB)
						    );
							 
ALU Alu (
													.Control(ALUControl),
													.A(SrcA),
													.B(SrcB),
													.Result(ALUResult)
        );
		  
Reg_param Result_register (
													.rst(reset), 
													.clk(clk), 
													.enable(1'b1), 
													.D(ALUResult), 
													.Q(ALUOut)
							);
							
							
Mux4x1 Result_mux (
								 .Selector(PCSrc),
								 .I_0(ALUResult),
								 .I_1(ALUOut),
								 //.I_2(ALUOut - 4),
								 .I_2(ALUOut),
								 .I_3(ALUResult - 4),
								 .Mux_Out(pc_next)
						   );
							
assign Op = op_q;
assign Funct3 = funct3_q;
assign Funct7 = funct7_q;
assign Zero = !ALUResult;

					
endmodule
